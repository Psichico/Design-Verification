package my_package;
import uvm_pkg::*;

`include "generate_sequence.sv"
`include "my_sequence.sv"
`include "sequencer.sv"
`include "driver.sv"
`include "monitor.sv"
`include "agent.sv"
`include "scoreboard.sv"
`include "my_environment.sv"
`include "test.sv"

endpackage
