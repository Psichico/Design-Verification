package my_package;
import uvm_pkg::*;

`include "/home/014512836/pal/273/monitor/generate_sequence.sv"
`include "/home/014512836/pal/273/monitor/my_sequence.sv"
`include "/home/014512836/pal/273/monitor/sequencer.sv"
`include "/home/014512836/pal/273/monitor/driver.sv"
`include "/home/014512836/pal/273/monitor/monitor.sv"
`include "/home/014512836/pal/273/monitor/monitor.sv"
`include "/home/014512836/pal/273/monitor/scoreboard.sv"
`include "/home/014512836/pal/273/monitor/my_environment.sv"
`include "/home/014512836/pal/273/monitor/test.sv"

endpackage
